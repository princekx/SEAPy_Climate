netcdf convert {  // CDL notation for a netCDF convert program

dimensions:         // dimension names and lengths are declared first
        lat = 64, lon = 129, level = 1, time = unlimited;

variables:          // variable types, names, shapes, attributes
        float   var(time,level,lat,lon);
                    var:long_name     = "variable";
        float     lat(lat), lon(lon), level(level);
                    lat:units       = "degrees";
                    lon:units       = "degrees";
        int   time(time);

data:                // optional data assignments
        level   = 1;
        lat     = -87.86, -85.10, -82.31, -79.53, -76.74, -73.95, -71.16,
                  -68.37, -65.58, -62.79, -60.00, -57.21, -54.42, -51.63, 
                  -48.84, -46.04, -43.25, -40.46, -37.67, -34.88, -32.09,
                  -29.30, -26.51, -23.72, -20.93, -18.14, -15.35, -12.56,
                   -9.77,  -6.98,  -4.19,  -1.40,   1.40,   4.19,   6.98,
                    9.77,  12.56,  15.35,  18.14,  20.93,  23.72,  26.51,
                   29.30,  32.09,  34.88,  37.67,  40.46,  43.25,  46.04,
                   48.84,  51.63,  54.42,  57.21,  60.00,  62.79,  65.58,
                   68.37,  71.16,  73.95,  76.74,  79.53,  82.31,  85.10,
                   87.86;
        lon     =   0.00,   2.81,   5.62,   8.44,  11.25,  14.06,  16.88,
                   19.69,  22.50,  25.31,  28.12,  30.94,  33.75,  36.56,
                   39.38,  42.19,  45.00,  47.81,  50.62,  53.44,  56.25,
                   59.06,  61.88,  64.69,  67.50,  70.31,  73.12,  75.94,
                   78.75,  81.56,  84.38,  87.19,  90.00,  92.81,  95.62,
                   98.44, 101.25, 104.06, 106.88, 109.69, 112.50, 115.31,
                  118.12, 120.94, 123.75, 126.56, 129.38, 132.19, 135.00,
                  137.81, 140.62, 143.44, 146.25, 149.06, 151.88, 154.69,
                  157.50, 160.31, 163.12, 165.94, 168.75, 171.56, 174.38,
                  177.19, 180.00, 182.81, 185.62, 188.44, 191.25, 194.06,
                  196.88, 199.69, 202.50, 205.31, 208.12, 210.94, 213.75,
                  216.56, 219.38, 222.19, 225.00, 227.81, 230.62, 233.44,
                  236.25, 239.06, 241.88, 244.69, 247.50, 250.31, 253.12,
                  255.94, 258.75, 261.56, 264.38, 267.19, 270.00, 272.81,
                  275.62, 278.44, 281.25, 284.06, 286.88, 289.69, 292.50,
                  295.31, 298.12, 300.94, 303.75, 306.56, 309.38, 312.19,
                  315.00, 317.81, 320.62, 323.44, 326.25, 329.06, 331.88,
                  334.69, 337.50, 340.31, 343.12, 345.94, 348.75, 351.56,
                  354.38, 357.19, 360.00;
        time    = 1,2,3,4,5,6,7;
}
